`timescale 1ns / 1ps

module VGA(
    input wire clk_25m,
    input wire clk_100m,
    input wire rst,
    input wire [31:0] pc,
    input wire [31:0] inst,
    input wire [31:0] alu_res,
    input wire mem_wen,
    input wire [31:0] dmem_o_data,
    input wire [31:0] dmem_i_data,
    input wire [31:0] dmem_addr,
    
    output wire hs,
    output wire vs,
    output wire [3:0] vga_r,
    output wire [3:0] vga_g,
    output wire [3:0] vga_b,

    input [32*32-1:0] regfile,
    input [31:0] alu_op1_val,
    input [31:0] alu_op2_val
    );
    wire [9:0] vga_x;
    wire [8:0] vga_y;
    wire video_on;
    VgaController vga_controller(
           .clk          (clk_25m      ),
           .rst          (rst          ),
           .vga_x        (vga_x        ),
           .vga_y        (vga_y        ),
           .hs           (hs           ),
           .vs           (vs           ),
           .video_on     (video_on     )
      );
 wire display_wen;
 wire [11:0] display_w_addr;
 wire [7:0] display_w_data;
 VgaDisplay vga_display(
          .clk          (clk_100m      ),
          .video_on     (video_on      ),
          .vga_x        (vga_x         ),
          .vga_y        (vga_y         ),
          .vga_r        (vga_r         ),
          .vga_g        (vga_g         ),
          .vga_b        (vga_b         ),
          .wen          (display_wen   ),
          .w_addr       (display_w_addr),
          .w_data       (display_w_data)
      );
 VgaDebugger vga_debugger(
         .clk           (clk_100m      ),
         .display_wen   (display_wen   ),
         .display_w_addr(display_w_addr),
         .display_w_data(display_w_data),
         .pc            (pc             ),
         .inst          (inst           ),
         .rs1           (               ),
         .rs1_val       (               ),
         .rs2           (               ),
         .rs2_val       (               ),
         .rd            (               ),
         .reg_i_data    (               ),
         .reg_wen       (               ),
         .is_imm        (               ),
         .is_auipc      (               ),
         .is_lui        (               ),
         .imm           (               ),
         .a_val         (alu_op1_val    ),
         .b_val         (alu_op2_val    ),
         .alu_ctrl      (               ),
         .cmp_ctrl      (               ),
         .alu_res       (alu_res        ),
         .cmp_res       (               ),
         .is_branch     (               ),
         .is_jal        (               ),
         .is_jalr       (               ),
         .do_branch     (               ),
         .pc_branch     (               ),
         .mem_wen       (mem_wen        ),
         .mem_ren       (               ),
         .dmem_o_data   (dmem_o_data    ),
         .dmem_i_data   (dmem_i_data    ),
         .dmem_addr     (dmem_addr      ),
         .csr_wen       (               ),
         .csr_ind       (               ),
         .csr_ctrl      (               ),
         .csr_r_data    (               ),
         .x0            (regfile[0*32+31 -: 32]),
         .ra            (regfile[1*32+31 -: 32]),
         .sp            (regfile[2*32+31 -: 32]),
         .gp            (regfile[3*32+31 -: 32]),
         .tp            (regfile[4*32+31 -: 32]),
         .t0            (regfile[5*32+31 -: 32]),
         .t1            (regfile[6*32+31 -: 32]),
         .t2            (regfile[7*32+31 -: 32]),
         .s0            (regfile[8*32+31 -: 32]),
         .s1            (regfile[9*32+31 -: 32]),
         .a0            (regfile[10*32+31 -: 32]),
         .a1            (regfile[11*32+31 -: 32]),
         .a2            (regfile[12*32+31 -: 32]),
         .a3            (regfile[13*32+31 -: 32]),
         .a4            (regfile[14*32+31 -: 32]),
         .a5            (regfile[15*32+31 -: 32]),
         .a6            (regfile[16*32+31 -: 32]),
         .a7            (regfile[17*32+31 -: 32]),
         .s2            (regfile[18*32+31 -: 32]),
         .s3            (regfile[19*32+31 -: 32]),
         .s4            (regfile[20*32+31 -: 32]),
         .s5            (regfile[21*32+31 -: 32]),
         .s6            (regfile[22*32+31 -: 32]),
         .s7            (regfile[23*32+31 -: 32]),
         .s8            (regfile[24*32+31 -: 32]),
         .s9            (regfile[25*32+31 -: 32]),
         .s10           (regfile[26*32+31 -: 32]),
         .s11           (regfile[27*32+31 -: 32]),
         .t3            (regfile[28*32+31 -: 32]),
         .t4            (regfile[29*32+31 -: 32]),
         .t5            (regfile[30*32+31 -: 32]),
         .t6            (regfile[31*32+31 -: 32]),
         .mstatus_o     (               ),
         .mcause_o      (               ),
         .mepc_o        (               ),
         .mtval_o       (               ),
         .mtvec_o       (               ),
         .mie_o         (               ),
         .mip_o         (               )
     );
endmodule

